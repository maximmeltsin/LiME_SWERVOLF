7c029073aaaa02b7
0000000000000067